//try after to implement at logic level. Or pipelined
module ALU (
    input logic [3:0] sel,
    input logic [3:0] A,
    input logic [3:0] B,
    input logic M,
    input logic Cn,
    output logic [3:0] F
);


